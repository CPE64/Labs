module 595SerialOuput(
  input     [8:0]     dataToSend,
  input               clk,

  output              serialOut,
  output              latch,
);

