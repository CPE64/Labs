//| This assertion will list an error if not met
assert (Logical statement)
    begin
    //<code-for-true-case>
    end
else
    begin
    //<code-for-false-case>
    end