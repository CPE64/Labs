  Adder #(
    .constant(SpecifiedConstant)
  )AdderDUT(
    .UserNumber(Number),
    .sum(Sum)
  );