  <Module>#(
    .<ParameterName>()
    )<InstanceName>(
    .<PortName>(<Wire>),
    .<PortName>(<Reg>)
  );