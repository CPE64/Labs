case(<StateRegister>)
    <Case 1>:<Statement>
    <Case 2>:<Statement>
    ....
    default:<Statement>