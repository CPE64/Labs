  //| This assertion will list an error if not met
  assert (Logical statement)
  <code-for-true-case>
  else
  <code-for-false-case>