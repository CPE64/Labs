  <Module><InstanceName>(
    .<PortName>(<Wire>),
    .<PortName>(<Reg>)
  );